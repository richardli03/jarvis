(
    show_hierarchy: None,
    show_menu: None,
    show_ticks: None,
    show_toolbar: None,
    show_tooltip: None,
    show_scope_tooltip: None,
    show_default_timeline: None,
    show_overview: None,
    show_statusbar: None,
    align_names_right: None,
    show_variable_indices: None,
    show_variable_direction: None,
    show_empty_scopes: None,
    show_parameters_in_scopes: None,
    highlight_focused: None,
    waves: Some((
        source: File("./sim_build/uart_main/uart_main.fst"),
        format: Fst,
        active_scope: Some(WaveScope((
            strs: [
                "uart_main",
            ],
        ))),
        items_tree: (
            items: [
                (
                    item_ref: (6),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (1),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (17),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (15),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (2),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (22),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (7),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (3),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (4),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (5),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (13),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (25),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (14),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (12),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (24),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (9),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (8),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (11),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (10),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (23),
                    level: 0,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (16),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (18),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (19),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
                (
                    item_ref: (20),
                    level: 1,
                    unfolded: true,
                    selected: false,
                ),
            ],
        ),
        displayed_items: {
            (22): Group((
                name: "receive",
                color: Some("Gray"),
                background_color: Some("Gray"),
                content: [],
                is_open: false,
            )),
            (16): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "tx",
                ),
                color: None,
                background_color: None,
                display_name: "tx",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (13): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_shift_en",
                ),
                color: None,
                background_color: None,
                display_name: "rx_shift_en",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (12): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_next_state",
                ),
                color: None,
                background_color: None,
                display_name: "rx_next_state [3:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (17): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "uart_clk",
                ),
                color: None,
                background_color: None,
                display_name: "uart_clk",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (4): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "read_ready",
                ),
                color: None,
                background_color: None,
                display_name: "read_ready",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (3): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "read_data",
                ),
                color: None,
                background_color: None,
                display_name: "read_data [7:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (6): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rst_n",
                ),
                color: None,
                background_color: None,
                display_name: "rst_n",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (20): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "write_valid",
                ),
                color: None,
                background_color: None,
                display_name: "write_valid",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (23): Group((
                name: "transmit",
                color: Some("Gray"),
                background_color: Some("Gray"),
                content: [],
                is_open: false,
            )),
            (24): Group((
                name: "receive_counters",
                color: Some("Gray"),
                background_color: Some("Gray"),
                content: [],
                is_open: false,
            )),
            (10): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_clk_counter",
                ),
                color: None,
                background_color: None,
                display_name: "rx_clk_counter [6:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (8): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_bit_counter",
                ),
                color: None,
                background_color: None,
                display_name: "rx_bit_counter [2:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (18): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "write_data",
                ),
                color: None,
                background_color: None,
                display_name: "write_data [7:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (25): Group((
                name: "receive_states",
                color: None,
                background_color: None,
                content: [],
                is_open: false,
            )),
            (9): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_bit_counter_rst_n",
                ),
                color: None,
                background_color: None,
                display_name: "rx_bit_counter_rst_n",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (14): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_state",
                ),
                color: None,
                background_color: None,
                display_name: "rx_state [3:0]",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (7): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx",
                ),
                color: None,
                background_color: None,
                display_name: "rx",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (2): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "mode",
                ),
                color: None,
                background_color: None,
                display_name: "mode",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (11): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "rx_clk_counter_rst_n",
                ),
                color: None,
                background_color: None,
                display_name: "rx_clk_counter_rst_n",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (15): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "sample_clk",
                ),
                color: None,
                background_color: None,
                display_name: "sample_clk",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (21): Group((
                name: "receive",
                color: None,
                background_color: None,
                content: [],
                is_open: false,
            )),
            (19): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "write_ready",
                ),
                color: None,
                background_color: None,
                display_name: "write_ready",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (1): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "clk",
                ),
                color: None,
                background_color: None,
                display_name: "clk",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
            (5): Variable((
                variable_ref: (
                    path: (
                        strs: [
                            "uart_main",
                        ],
                    ),
                    name: "read_valid",
                ),
                color: None,
                background_color: None,
                display_name: "read_valid",
                display_name_type: Unique,
                manual_name: None,
                format: None,
                field_formats: [],
            )),
        },
        display_item_ref_counter: 25,
        viewports: [
            (
                curr_left: (0.0),
                curr_right: (1.3999999999999997),
                target_left: (0.0),
                target_right: (1.0),
                move_start_left: (0.0),
                move_start_right: (1.0),
                move_duration: None,
                move_strategy: Instant,
            ),
        ],
        cursor: Some((1, [
            295107,
        ])),
        markers: {},
        focused_item: None,
        focused_transaction: (None, None),
        default_variable_name_type: Unique,
        scroll_offset: 0.0,
        display_variable_indices: true,
        graphics: {},
    )),
    drag_started: false,
    drag_source_idx: None,
    drag_target_idx: Some((
        before: (10),
        level: 1,
    )),
    previous_waves: None,
    count: None,
    blacklisted_translators: [],
    show_about: false,
    show_keys: false,
    show_gestures: false,
    show_quick_start: false,
    show_license: false,
    show_performance: false,
    show_logs: false,
    show_cursor_window: false,
    wanted_timeunit: PicoSeconds,
    time_string_format: None,
    show_url_entry: false,
    variable_name_filter_focused: false,
    variable_name_filter_type: Fuzzy,
    variable_name_filter_case_insensitive: true,
    rename_target: None,
    sidepanel_width: Some(297.96875),
    ui_zoom_factor: None,
)